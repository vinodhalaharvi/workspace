entity mac_test is

end entity mac_test;
