test_bench-join.vhdl