entity to_fp_test is

end entity to_fp_test;
