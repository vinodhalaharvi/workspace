package pk_04_02 is

  subtype halfword is bit_vector(0 to 15);

end package pk_04_02;
