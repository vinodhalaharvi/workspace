join.vhdl