fork.vhdl