queue.vhdl