server.vhdl