test_bench-join_synth.vhdl