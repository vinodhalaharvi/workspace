entity test_bench is

end entity test_bench;
