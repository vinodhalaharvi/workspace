random.vhdl