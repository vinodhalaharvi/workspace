test_bench-source.vhdl