server-behavior.vhdl