entity disk_system is

end entity disk_system;

