waiting_token_fifo_adt.vhdl