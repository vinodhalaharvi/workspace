source.vhdl