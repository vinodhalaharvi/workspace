test_bench-fork.vhdl