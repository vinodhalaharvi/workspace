disk_system-queue_net.vhdl