package pk_04_01 is

  subtype coeff_ram_address is integer range 0 to 63;

end package pk_04_01;
