queue-behavior.vhdl