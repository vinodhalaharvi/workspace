token_fifo_adt-body.vhdl