source-behavior.vhdl