test_bench-queue_server.vhdl