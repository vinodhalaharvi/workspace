test_bench-sink.vhdl