test_bench.vhdl