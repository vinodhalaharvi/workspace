package test_bench_03_02 is

  -- following type used in Figure 3-02

  -- code from book:

  type sel_range is range 0 to 3;

  -- end of code from book

end package test_bench_03_02;
