fork-behavior.vhdl