disk_system.vhdl