-- not in book

use work.tb_05_13.all;

-- end not in book

entity adder is
  port ( a : in word;
         b : in word;
         sum : out word );
end entity adder;
