entity computer is

end entity computer;
