sink.vhdl