qsim_types.vhdl