queue_types.vhdl