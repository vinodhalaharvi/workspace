random-body.vhdl