sink-behavior.vhdl