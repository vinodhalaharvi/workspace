token_fifo_adt.vhdl