join-behavior.vhdl