qsim_types-body.vhdl